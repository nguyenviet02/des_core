VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO des_core
  CLASS BLOCK ;
  FOREIGN des_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 1200.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.740 10.640 640.340 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 792.340 10.640 793.940 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 945.940 10.640 947.540 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1099.540 10.640 1101.140 1188.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 1194.400 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 1194.400 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 1194.400 337.990 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 489.570 1194.400 491.170 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 642.750 1194.400 644.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 795.930 1194.400 797.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 949.110 1194.400 950.710 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1102.290 1194.400 1103.890 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1188.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 1194.400 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 1194.400 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 1194.400 334.690 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 486.270 1194.400 487.870 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 639.450 1194.400 641.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 792.630 1194.400 794.230 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 945.810 1194.400 947.410 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1098.990 1194.400 1100.590 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END clk
  PIN des_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 438.640 1200.000 439.240 ;
    END
  END des_data[0]
  PIN des_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END des_data[10]
  PIN des_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END des_data[11]
  PIN des_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 592.570 1196.000 592.850 1200.000 ;
    END
  END des_data[12]
  PIN des_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END des_data[13]
  PIN des_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END des_data[14]
  PIN des_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.840 4.000 772.440 ;
    END
  END des_data[15]
  PIN des_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 705.270 1196.000 705.550 1200.000 ;
    END
  END des_data[16]
  PIN des_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 595.790 1196.000 596.070 1200.000 ;
    END
  END des_data[17]
  PIN des_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 452.240 1200.000 452.840 ;
    END
  END des_data[18]
  PIN des_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 527.040 1200.000 527.640 ;
    END
  END des_data[19]
  PIN des_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 476.040 1200.000 476.640 ;
    END
  END des_data[1]
  PIN des_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END des_data[20]
  PIN des_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END des_data[21]
  PIN des_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END des_data[22]
  PIN des_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END des_data[23]
  PIN des_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 599.010 1196.000 599.290 1200.000 ;
    END
  END des_data[24]
  PIN des_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 679.510 1196.000 679.790 1200.000 ;
    END
  END des_data[25]
  PIN des_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 601.840 1200.000 602.440 ;
    END
  END des_data[26]
  PIN des_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 510.040 1200.000 510.640 ;
    END
  END des_data[27]
  PIN des_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 685.950 1196.000 686.230 1200.000 ;
    END
  END des_data[28]
  PIN des_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END des_data[29]
  PIN des_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END des_data[2]
  PIN des_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 521.730 0.000 522.010 4.000 ;
    END
  END des_data[30]
  PIN des_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END des_data[31]
  PIN des_data[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 472.640 1200.000 473.240 ;
    END
  END des_data[32]
  PIN des_data[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 479.440 1200.000 480.040 ;
    END
  END des_data[33]
  PIN des_data[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 530.440 1200.000 531.040 ;
    END
  END des_data[34]
  PIN des_data[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 442.040 1200.000 442.640 ;
    END
  END des_data[35]
  PIN des_data[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END des_data[36]
  PIN des_data[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END des_data[37]
  PIN des_data[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 660.190 1196.000 660.470 1200.000 ;
    END
  END des_data[38]
  PIN des_data[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 634.430 1196.000 634.710 1200.000 ;
    END
  END des_data[39]
  PIN des_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END des_data[3]
  PIN des_data[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 669.850 1196.000 670.130 1200.000 ;
    END
  END des_data[40]
  PIN des_data[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 676.290 1196.000 676.570 1200.000 ;
    END
  END des_data[41]
  PIN des_data[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 493.040 1200.000 493.640 ;
    END
  END des_data[42]
  PIN des_data[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 482.840 1200.000 483.440 ;
    END
  END des_data[43]
  PIN des_data[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END des_data[44]
  PIN des_data[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.840 4.000 602.440 ;
    END
  END des_data[45]
  PIN des_data[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END des_data[46]
  PIN des_data[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END des_data[47]
  PIN des_data[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 624.770 1196.000 625.050 1200.000 ;
    END
  END des_data[48]
  PIN des_data[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 666.630 1196.000 666.910 1200.000 ;
    END
  END des_data[49]
  PIN des_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END des_data[4]
  PIN des_data[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END des_data[50]
  PIN des_data[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 506.640 1200.000 507.240 ;
    END
  END des_data[51]
  PIN des_data[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 695.610 1196.000 695.890 1200.000 ;
    END
  END des_data[52]
  PIN des_data[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 608.670 1196.000 608.950 1200.000 ;
    END
  END des_data[53]
  PIN des_data[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END des_data[54]
  PIN des_data[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END des_data[55]
  PIN des_data[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 731.030 1196.000 731.310 1200.000 ;
    END
  END des_data[56]
  PIN des_data[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 714.930 1196.000 715.210 1200.000 ;
    END
  END des_data[57]
  PIN des_data[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 611.890 1196.000 612.170 1200.000 ;
    END
  END des_data[58]
  PIN des_data[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 537.240 1200.000 537.840 ;
    END
  END des_data[59]
  PIN des_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END des_data[5]
  PIN des_data[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END des_data[60]
  PIN des_data[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 676.640 4.000 677.240 ;
    END
  END des_data[61]
  PIN des_data[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END des_data[62]
  PIN des_data[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END des_data[63]
  PIN des_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 627.990 1196.000 628.270 1200.000 ;
    END
  END des_data[6]
  PIN des_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 631.210 1196.000 631.490 1200.000 ;
    END
  END des_data[7]
  PIN des_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 708.490 1196.000 708.770 1200.000 ;
    END
  END des_data[8]
  PIN des_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 724.590 1196.000 724.870 1200.000 ;
    END
  END des_data[9]
  PIN des_decipher_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END des_decipher_en
  PIN des_encipher_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END des_encipher_en
  PIN des_key_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END des_key_in[0]
  PIN des_key_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 608.640 1200.000 609.240 ;
    END
  END des_key_in[10]
  PIN des_key_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 571.240 1200.000 571.840 ;
    END
  END des_key_in[11]
  PIN des_key_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 615.440 4.000 616.040 ;
    END
  END des_key_in[12]
  PIN des_key_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END des_key_in[13]
  PIN des_key_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END des_key_in[14]
  PIN des_key_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END des_key_in[15]
  PIN des_key_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END des_key_in[16]
  PIN des_key_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 561.040 1200.000 561.640 ;
    END
  END des_key_in[17]
  PIN des_key_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 605.240 1200.000 605.840 ;
    END
  END des_key_in[18]
  PIN des_key_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 516.840 1200.000 517.440 ;
    END
  END des_key_in[19]
  PIN des_key_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 598.440 1200.000 599.040 ;
    END
  END des_key_in[1]
  PIN des_key_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END des_key_in[20]
  PIN des_key_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 710.640 4.000 711.240 ;
    END
  END des_key_in[21]
  PIN des_key_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 683.440 4.000 684.040 ;
    END
  END des_key_in[22]
  PIN des_key_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END des_key_in[23]
  PIN des_key_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END des_key_in[24]
  PIN des_key_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 647.310 1196.000 647.590 1200.000 ;
    END
  END des_key_in[25]
  PIN des_key_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 544.040 1200.000 544.640 ;
    END
  END des_key_in[26]
  PIN des_key_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 496.440 1200.000 497.040 ;
    END
  END des_key_in[27]
  PIN des_key_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END des_key_in[28]
  PIN des_key_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END des_key_in[29]
  PIN des_key_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 567.840 1200.000 568.440 ;
    END
  END des_key_in[2]
  PIN des_key_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.840 4.000 704.440 ;
    END
  END des_key_in[30]
  PIN des_key_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END des_key_in[31]
  PIN des_key_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END des_key_in[32]
  PIN des_key_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 564.440 1200.000 565.040 ;
    END
  END des_key_in[33]
  PIN des_key_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 574.640 1200.000 575.240 ;
    END
  END des_key_in[34]
  PIN des_key_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 513.440 1200.000 514.040 ;
    END
  END des_key_in[35]
  PIN des_key_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 547.440 1200.000 548.040 ;
    END
  END des_key_in[36]
  PIN des_key_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END des_key_in[37]
  PIN des_key_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END des_key_in[38]
  PIN des_key_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END des_key_in[39]
  PIN des_key_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 520.240 1200.000 520.840 ;
    END
  END des_key_in[3]
  PIN des_key_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END des_key_in[40]
  PIN des_key_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 682.730 1196.000 683.010 1200.000 ;
    END
  END des_key_in[41]
  PIN des_key_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 588.240 1200.000 588.840 ;
    END
  END des_key_in[42]
  PIN des_key_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 581.440 1200.000 582.040 ;
    END
  END des_key_in[43]
  PIN des_key_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 540.640 1200.000 541.240 ;
    END
  END des_key_in[44]
  PIN des_key_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.040 4.000 629.640 ;
    END
  END des_key_in[45]
  PIN des_key_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.240 4.000 656.840 ;
    END
  END des_key_in[46]
  PIN des_key_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END des_key_in[47]
  PIN des_key_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END des_key_in[48]
  PIN des_key_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 595.040 1200.000 595.640 ;
    END
  END des_key_in[49]
  PIN des_key_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END des_key_in[4]
  PIN des_key_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 554.240 1200.000 554.840 ;
    END
  END des_key_in[50]
  PIN des_key_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 499.840 1200.000 500.440 ;
    END
  END des_key_in[51]
  PIN des_key_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 533.840 1200.000 534.440 ;
    END
  END des_key_in[52]
  PIN des_key_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END des_key_in[53]
  PIN des_key_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 649.440 4.000 650.040 ;
    END
  END des_key_in[54]
  PIN des_key_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.240 4.000 690.840 ;
    END
  END des_key_in[55]
  PIN des_key_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END des_key_in[56]
  PIN des_key_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 689.170 1196.000 689.450 1200.000 ;
    END
  END des_key_in[57]
  PIN des_key_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 550.840 1200.000 551.440 ;
    END
  END des_key_in[58]
  PIN des_key_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 523.640 1200.000 524.240 ;
    END
  END des_key_in[59]
  PIN des_key_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END des_key_in[5]
  PIN des_key_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 591.640 1200.000 592.240 ;
    END
  END des_key_in[60]
  PIN des_key_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 608.640 4.000 609.240 ;
    END
  END des_key_in[61]
  PIN des_key_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END des_key_in[62]
  PIN des_key_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END des_key_in[63]
  PIN des_key_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END des_key_in[6]
  PIN des_key_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 505.630 0.000 505.910 4.000 ;
    END
  END des_key_in[7]
  PIN des_key_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END des_key_in[8]
  PIN des_key_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 557.640 1200.000 558.240 ;
    END
  END des_key_in[9]
  PIN desc_ready
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END desc_ready
  PIN desc_result[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 462.440 1200.000 463.040 ;
    END
  END desc_result[0]
  PIN desc_result[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 4.000 ;
    END
  END desc_result[10]
  PIN desc_result[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END desc_result[11]
  PIN desc_result[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 751.440 4.000 752.040 ;
    END
  END desc_result[12]
  PIN desc_result[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 744.640 4.000 745.240 ;
    END
  END desc_result[13]
  PIN desc_result[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END desc_result[14]
  PIN desc_result[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.840 4.000 670.440 ;
    END
  END desc_result[15]
  PIN desc_result[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 702.050 1196.000 702.330 1200.000 ;
    END
  END desc_result[16]
  PIN desc_result[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 711.710 1196.000 711.990 1200.000 ;
    END
  END desc_result[17]
  PIN desc_result[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 455.640 1200.000 456.240 ;
    END
  END desc_result[18]
  PIN desc_result[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 459.040 1200.000 459.640 ;
    END
  END desc_result[19]
  PIN desc_result[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 469.240 1200.000 469.840 ;
    END
  END desc_result[1]
  PIN desc_result[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END desc_result[20]
  PIN desc_result[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.240 4.000 622.840 ;
    END
  END desc_result[21]
  PIN desc_result[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END desc_result[22]
  PIN desc_result[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END desc_result[23]
  PIN desc_result[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 621.550 1196.000 621.830 1200.000 ;
    END
  END desc_result[24]
  PIN desc_result[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 637.650 1196.000 637.930 1200.000 ;
    END
  END desc_result[25]
  PIN desc_result[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 584.840 1200.000 585.440 ;
    END
  END desc_result[26]
  PIN desc_result[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 578.040 1200.000 578.640 ;
    END
  END desc_result[27]
  PIN desc_result[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 650.530 1196.000 650.810 1200.000 ;
    END
  END desc_result[28]
  PIN desc_result[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 656.970 1196.000 657.250 1200.000 ;
    END
  END desc_result[29]
  PIN desc_result[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END desc_result[2]
  PIN desc_result[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END desc_result[30]
  PIN desc_result[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END desc_result[31]
  PIN desc_result[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 465.840 1200.000 466.440 ;
    END
  END desc_result[32]
  PIN desc_result[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 448.840 1200.000 449.440 ;
    END
  END desc_result[33]
  PIN desc_result[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 445.440 1200.000 446.040 ;
    END
  END desc_result[34]
  PIN desc_result[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 503.240 1200.000 503.840 ;
    END
  END desc_result[35]
  PIN desc_result[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END desc_result[36]
  PIN desc_result[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END desc_result[37]
  PIN desc_result[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 653.750 1196.000 654.030 1200.000 ;
    END
  END desc_result[38]
  PIN desc_result[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 644.090 1196.000 644.370 1200.000 ;
    END
  END desc_result[39]
  PIN desc_result[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 4.000 ;
    END
  END desc_result[3]
  PIN desc_result[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 673.070 1196.000 673.350 1200.000 ;
    END
  END desc_result[40]
  PIN desc_result[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 698.830 1196.000 699.110 1200.000 ;
    END
  END desc_result[41]
  PIN desc_result[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 489.640 1200.000 490.240 ;
    END
  END desc_result[42]
  PIN desc_result[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 486.240 1200.000 486.840 ;
    END
  END desc_result[43]
  PIN desc_result[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END desc_result[44]
  PIN desc_result[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END desc_result[45]
  PIN desc_result[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END desc_result[46]
  PIN desc_result[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END desc_result[47]
  PIN desc_result[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 602.230 1196.000 602.510 1200.000 ;
    END
  END desc_result[48]
  PIN desc_result[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 605.450 1196.000 605.730 1200.000 ;
    END
  END desc_result[49]
  PIN desc_result[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END desc_result[4]
  PIN desc_result[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END desc_result[50]
  PIN desc_result[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END desc_result[51]
  PIN desc_result[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 663.410 1196.000 663.690 1200.000 ;
    END
  END desc_result[52]
  PIN desc_result[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 692.390 1196.000 692.670 1200.000 ;
    END
  END desc_result[53]
  PIN desc_result[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END desc_result[54]
  PIN desc_result[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END desc_result[55]
  PIN desc_result[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 734.250 1196.000 734.530 1200.000 ;
    END
  END desc_result[56]
  PIN desc_result[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 727.810 1196.000 728.090 1200.000 ;
    END
  END desc_result[57]
  PIN desc_result[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 612.040 1200.000 612.640 ;
    END
  END desc_result[58]
  PIN desc_result[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 615.110 1196.000 615.390 1200.000 ;
    END
  END desc_result[59]
  PIN desc_result[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.240 4.000 724.840 ;
    END
  END desc_result[5]
  PIN desc_result[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END desc_result[60]
  PIN desc_result[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END desc_result[61]
  PIN desc_result[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END desc_result[62]
  PIN desc_result[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END desc_result[63]
  PIN desc_result[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 640.870 1196.000 641.150 1200.000 ;
    END
  END desc_result[6]
  PIN desc_result[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 618.330 1196.000 618.610 1200.000 ;
    END
  END desc_result[7]
  PIN desc_result[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 718.150 1196.000 718.430 1200.000 ;
    END
  END desc_result[8]
  PIN desc_result[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 721.370 1196.000 721.650 1200.000 ;
    END
  END desc_result[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 486.310 0.000 486.590 4.000 ;
    END
  END rst_n
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1194.160 1188.725 ;
      LAYER met1 ;
        RECT 4.210 10.640 1194.160 1189.960 ;
      LAYER met2 ;
        RECT 4.230 1195.720 592.290 1196.530 ;
        RECT 593.130 1195.720 595.510 1196.530 ;
        RECT 596.350 1195.720 598.730 1196.530 ;
        RECT 599.570 1195.720 601.950 1196.530 ;
        RECT 602.790 1195.720 605.170 1196.530 ;
        RECT 606.010 1195.720 608.390 1196.530 ;
        RECT 609.230 1195.720 611.610 1196.530 ;
        RECT 612.450 1195.720 614.830 1196.530 ;
        RECT 615.670 1195.720 618.050 1196.530 ;
        RECT 618.890 1195.720 621.270 1196.530 ;
        RECT 622.110 1195.720 624.490 1196.530 ;
        RECT 625.330 1195.720 627.710 1196.530 ;
        RECT 628.550 1195.720 630.930 1196.530 ;
        RECT 631.770 1195.720 634.150 1196.530 ;
        RECT 634.990 1195.720 637.370 1196.530 ;
        RECT 638.210 1195.720 640.590 1196.530 ;
        RECT 641.430 1195.720 643.810 1196.530 ;
        RECT 644.650 1195.720 647.030 1196.530 ;
        RECT 647.870 1195.720 650.250 1196.530 ;
        RECT 651.090 1195.720 653.470 1196.530 ;
        RECT 654.310 1195.720 656.690 1196.530 ;
        RECT 657.530 1195.720 659.910 1196.530 ;
        RECT 660.750 1195.720 663.130 1196.530 ;
        RECT 663.970 1195.720 666.350 1196.530 ;
        RECT 667.190 1195.720 669.570 1196.530 ;
        RECT 670.410 1195.720 672.790 1196.530 ;
        RECT 673.630 1195.720 676.010 1196.530 ;
        RECT 676.850 1195.720 679.230 1196.530 ;
        RECT 680.070 1195.720 682.450 1196.530 ;
        RECT 683.290 1195.720 685.670 1196.530 ;
        RECT 686.510 1195.720 688.890 1196.530 ;
        RECT 689.730 1195.720 692.110 1196.530 ;
        RECT 692.950 1195.720 695.330 1196.530 ;
        RECT 696.170 1195.720 698.550 1196.530 ;
        RECT 699.390 1195.720 701.770 1196.530 ;
        RECT 702.610 1195.720 704.990 1196.530 ;
        RECT 705.830 1195.720 708.210 1196.530 ;
        RECT 709.050 1195.720 711.430 1196.530 ;
        RECT 712.270 1195.720 714.650 1196.530 ;
        RECT 715.490 1195.720 717.870 1196.530 ;
        RECT 718.710 1195.720 721.090 1196.530 ;
        RECT 721.930 1195.720 724.310 1196.530 ;
        RECT 725.150 1195.720 727.530 1196.530 ;
        RECT 728.370 1195.720 730.750 1196.530 ;
        RECT 731.590 1195.720 733.970 1196.530 ;
        RECT 734.810 1195.720 1192.690 1196.530 ;
        RECT 4.230 4.280 1192.690 1195.720 ;
        RECT 4.230 3.670 6.250 4.280 ;
        RECT 7.090 3.670 9.470 4.280 ;
        RECT 10.310 3.670 12.690 4.280 ;
        RECT 13.530 3.670 15.910 4.280 ;
        RECT 16.750 3.670 19.130 4.280 ;
        RECT 19.970 3.670 22.350 4.280 ;
        RECT 23.190 3.670 453.830 4.280 ;
        RECT 454.670 3.670 457.050 4.280 ;
        RECT 457.890 3.670 460.270 4.280 ;
        RECT 461.110 3.670 463.490 4.280 ;
        RECT 464.330 3.670 466.710 4.280 ;
        RECT 467.550 3.670 469.930 4.280 ;
        RECT 470.770 3.670 473.150 4.280 ;
        RECT 473.990 3.670 476.370 4.280 ;
        RECT 477.210 3.670 479.590 4.280 ;
        RECT 480.430 3.670 482.810 4.280 ;
        RECT 483.650 3.670 486.030 4.280 ;
        RECT 486.870 3.670 492.470 4.280 ;
        RECT 493.310 3.670 495.690 4.280 ;
        RECT 496.530 3.670 498.910 4.280 ;
        RECT 499.750 3.670 502.130 4.280 ;
        RECT 502.970 3.670 505.350 4.280 ;
        RECT 506.190 3.670 508.570 4.280 ;
        RECT 509.410 3.670 511.790 4.280 ;
        RECT 512.630 3.670 515.010 4.280 ;
        RECT 515.850 3.670 518.230 4.280 ;
        RECT 519.070 3.670 521.450 4.280 ;
        RECT 522.290 3.670 524.670 4.280 ;
        RECT 525.510 3.670 527.890 4.280 ;
        RECT 528.730 3.670 531.110 4.280 ;
        RECT 531.950 3.670 534.330 4.280 ;
        RECT 535.170 3.670 537.550 4.280 ;
        RECT 538.390 3.670 540.770 4.280 ;
        RECT 541.610 3.670 543.990 4.280 ;
        RECT 544.830 3.670 547.210 4.280 ;
        RECT 548.050 3.670 550.430 4.280 ;
        RECT 551.270 3.670 553.650 4.280 ;
        RECT 554.490 3.670 556.870 4.280 ;
        RECT 557.710 3.670 560.090 4.280 ;
        RECT 560.930 3.670 563.310 4.280 ;
        RECT 564.150 3.670 566.530 4.280 ;
        RECT 567.370 3.670 576.190 4.280 ;
        RECT 577.030 3.670 579.410 4.280 ;
        RECT 580.250 3.670 582.630 4.280 ;
        RECT 583.470 3.670 1192.690 4.280 ;
      LAYER met3 ;
        RECT 3.990 772.840 1196.000 1188.805 ;
        RECT 4.400 771.440 1196.000 772.840 ;
        RECT 3.990 769.440 1196.000 771.440 ;
        RECT 4.400 768.040 1196.000 769.440 ;
        RECT 3.990 766.040 1196.000 768.040 ;
        RECT 4.400 764.640 1196.000 766.040 ;
        RECT 3.990 762.640 1196.000 764.640 ;
        RECT 4.400 761.240 1196.000 762.640 ;
        RECT 3.990 759.240 1196.000 761.240 ;
        RECT 4.400 757.840 1196.000 759.240 ;
        RECT 3.990 755.840 1196.000 757.840 ;
        RECT 4.400 754.440 1196.000 755.840 ;
        RECT 3.990 752.440 1196.000 754.440 ;
        RECT 4.400 751.040 1196.000 752.440 ;
        RECT 3.990 749.040 1196.000 751.040 ;
        RECT 4.400 747.640 1196.000 749.040 ;
        RECT 3.990 745.640 1196.000 747.640 ;
        RECT 4.400 744.240 1196.000 745.640 ;
        RECT 3.990 742.240 1196.000 744.240 ;
        RECT 4.400 740.840 1196.000 742.240 ;
        RECT 3.990 738.840 1196.000 740.840 ;
        RECT 4.400 737.440 1196.000 738.840 ;
        RECT 3.990 735.440 1196.000 737.440 ;
        RECT 4.400 734.040 1196.000 735.440 ;
        RECT 3.990 732.040 1196.000 734.040 ;
        RECT 4.400 730.640 1196.000 732.040 ;
        RECT 3.990 728.640 1196.000 730.640 ;
        RECT 4.400 727.240 1196.000 728.640 ;
        RECT 3.990 725.240 1196.000 727.240 ;
        RECT 4.400 723.840 1196.000 725.240 ;
        RECT 3.990 721.840 1196.000 723.840 ;
        RECT 4.400 720.440 1196.000 721.840 ;
        RECT 3.990 718.440 1196.000 720.440 ;
        RECT 4.400 717.040 1196.000 718.440 ;
        RECT 3.990 715.040 1196.000 717.040 ;
        RECT 4.400 713.640 1196.000 715.040 ;
        RECT 3.990 711.640 1196.000 713.640 ;
        RECT 4.400 710.240 1196.000 711.640 ;
        RECT 3.990 708.240 1196.000 710.240 ;
        RECT 4.400 706.840 1196.000 708.240 ;
        RECT 3.990 704.840 1196.000 706.840 ;
        RECT 4.400 703.440 1196.000 704.840 ;
        RECT 3.990 701.440 1196.000 703.440 ;
        RECT 4.400 700.040 1196.000 701.440 ;
        RECT 3.990 698.040 1196.000 700.040 ;
        RECT 4.400 696.640 1196.000 698.040 ;
        RECT 3.990 694.640 1196.000 696.640 ;
        RECT 4.400 693.240 1196.000 694.640 ;
        RECT 3.990 691.240 1196.000 693.240 ;
        RECT 4.400 689.840 1196.000 691.240 ;
        RECT 3.990 687.840 1196.000 689.840 ;
        RECT 4.400 686.440 1196.000 687.840 ;
        RECT 3.990 684.440 1196.000 686.440 ;
        RECT 4.400 683.040 1196.000 684.440 ;
        RECT 3.990 681.040 1196.000 683.040 ;
        RECT 4.400 679.640 1196.000 681.040 ;
        RECT 3.990 677.640 1196.000 679.640 ;
        RECT 4.400 676.240 1196.000 677.640 ;
        RECT 3.990 674.240 1196.000 676.240 ;
        RECT 4.400 672.840 1196.000 674.240 ;
        RECT 3.990 670.840 1196.000 672.840 ;
        RECT 4.400 669.440 1196.000 670.840 ;
        RECT 3.990 667.440 1196.000 669.440 ;
        RECT 4.400 666.040 1196.000 667.440 ;
        RECT 3.990 664.040 1196.000 666.040 ;
        RECT 4.400 662.640 1196.000 664.040 ;
        RECT 3.990 660.640 1196.000 662.640 ;
        RECT 4.400 659.240 1196.000 660.640 ;
        RECT 3.990 657.240 1196.000 659.240 ;
        RECT 4.400 655.840 1196.000 657.240 ;
        RECT 3.990 653.840 1196.000 655.840 ;
        RECT 4.400 652.440 1196.000 653.840 ;
        RECT 3.990 650.440 1196.000 652.440 ;
        RECT 4.400 649.040 1196.000 650.440 ;
        RECT 3.990 647.040 1196.000 649.040 ;
        RECT 4.400 645.640 1196.000 647.040 ;
        RECT 3.990 643.640 1196.000 645.640 ;
        RECT 4.400 642.240 1196.000 643.640 ;
        RECT 3.990 640.240 1196.000 642.240 ;
        RECT 4.400 638.840 1196.000 640.240 ;
        RECT 3.990 636.840 1196.000 638.840 ;
        RECT 4.400 635.440 1196.000 636.840 ;
        RECT 3.990 633.440 1196.000 635.440 ;
        RECT 4.400 632.040 1196.000 633.440 ;
        RECT 3.990 630.040 1196.000 632.040 ;
        RECT 4.400 628.640 1196.000 630.040 ;
        RECT 3.990 626.640 1196.000 628.640 ;
        RECT 4.400 625.240 1196.000 626.640 ;
        RECT 3.990 623.240 1196.000 625.240 ;
        RECT 4.400 621.840 1196.000 623.240 ;
        RECT 3.990 619.840 1196.000 621.840 ;
        RECT 4.400 618.440 1196.000 619.840 ;
        RECT 3.990 616.440 1196.000 618.440 ;
        RECT 4.400 615.040 1196.000 616.440 ;
        RECT 3.990 613.040 1196.000 615.040 ;
        RECT 4.400 611.640 1195.600 613.040 ;
        RECT 3.990 609.640 1196.000 611.640 ;
        RECT 4.400 608.240 1195.600 609.640 ;
        RECT 3.990 606.240 1196.000 608.240 ;
        RECT 4.400 604.840 1195.600 606.240 ;
        RECT 3.990 602.840 1196.000 604.840 ;
        RECT 4.400 601.440 1195.600 602.840 ;
        RECT 3.990 599.440 1196.000 601.440 ;
        RECT 4.400 598.040 1195.600 599.440 ;
        RECT 3.990 596.040 1196.000 598.040 ;
        RECT 4.400 594.640 1195.600 596.040 ;
        RECT 3.990 592.640 1196.000 594.640 ;
        RECT 4.400 591.240 1195.600 592.640 ;
        RECT 3.990 589.240 1196.000 591.240 ;
        RECT 3.990 587.840 1195.600 589.240 ;
        RECT 3.990 585.840 1196.000 587.840 ;
        RECT 3.990 584.440 1195.600 585.840 ;
        RECT 3.990 582.440 1196.000 584.440 ;
        RECT 3.990 581.040 1195.600 582.440 ;
        RECT 3.990 579.040 1196.000 581.040 ;
        RECT 3.990 577.640 1195.600 579.040 ;
        RECT 3.990 575.640 1196.000 577.640 ;
        RECT 3.990 574.240 1195.600 575.640 ;
        RECT 3.990 572.240 1196.000 574.240 ;
        RECT 3.990 570.840 1195.600 572.240 ;
        RECT 3.990 568.840 1196.000 570.840 ;
        RECT 3.990 567.440 1195.600 568.840 ;
        RECT 3.990 565.440 1196.000 567.440 ;
        RECT 3.990 564.040 1195.600 565.440 ;
        RECT 3.990 562.040 1196.000 564.040 ;
        RECT 3.990 560.640 1195.600 562.040 ;
        RECT 3.990 558.640 1196.000 560.640 ;
        RECT 3.990 557.240 1195.600 558.640 ;
        RECT 3.990 555.240 1196.000 557.240 ;
        RECT 3.990 553.840 1195.600 555.240 ;
        RECT 3.990 551.840 1196.000 553.840 ;
        RECT 3.990 550.440 1195.600 551.840 ;
        RECT 3.990 548.440 1196.000 550.440 ;
        RECT 3.990 547.040 1195.600 548.440 ;
        RECT 3.990 545.040 1196.000 547.040 ;
        RECT 3.990 543.640 1195.600 545.040 ;
        RECT 3.990 541.640 1196.000 543.640 ;
        RECT 3.990 540.240 1195.600 541.640 ;
        RECT 3.990 538.240 1196.000 540.240 ;
        RECT 3.990 536.840 1195.600 538.240 ;
        RECT 3.990 534.840 1196.000 536.840 ;
        RECT 3.990 533.440 1195.600 534.840 ;
        RECT 3.990 531.440 1196.000 533.440 ;
        RECT 3.990 530.040 1195.600 531.440 ;
        RECT 3.990 528.040 1196.000 530.040 ;
        RECT 3.990 526.640 1195.600 528.040 ;
        RECT 3.990 524.640 1196.000 526.640 ;
        RECT 3.990 523.240 1195.600 524.640 ;
        RECT 3.990 521.240 1196.000 523.240 ;
        RECT 3.990 519.840 1195.600 521.240 ;
        RECT 3.990 517.840 1196.000 519.840 ;
        RECT 3.990 516.440 1195.600 517.840 ;
        RECT 3.990 514.440 1196.000 516.440 ;
        RECT 3.990 513.040 1195.600 514.440 ;
        RECT 3.990 511.040 1196.000 513.040 ;
        RECT 3.990 509.640 1195.600 511.040 ;
        RECT 3.990 507.640 1196.000 509.640 ;
        RECT 3.990 506.240 1195.600 507.640 ;
        RECT 3.990 504.240 1196.000 506.240 ;
        RECT 3.990 502.840 1195.600 504.240 ;
        RECT 3.990 500.840 1196.000 502.840 ;
        RECT 3.990 499.440 1195.600 500.840 ;
        RECT 3.990 497.440 1196.000 499.440 ;
        RECT 3.990 496.040 1195.600 497.440 ;
        RECT 3.990 494.040 1196.000 496.040 ;
        RECT 3.990 492.640 1195.600 494.040 ;
        RECT 3.990 490.640 1196.000 492.640 ;
        RECT 3.990 489.240 1195.600 490.640 ;
        RECT 3.990 487.240 1196.000 489.240 ;
        RECT 3.990 485.840 1195.600 487.240 ;
        RECT 3.990 483.840 1196.000 485.840 ;
        RECT 3.990 482.440 1195.600 483.840 ;
        RECT 3.990 480.440 1196.000 482.440 ;
        RECT 3.990 479.040 1195.600 480.440 ;
        RECT 3.990 477.040 1196.000 479.040 ;
        RECT 3.990 475.640 1195.600 477.040 ;
        RECT 3.990 473.640 1196.000 475.640 ;
        RECT 3.990 472.240 1195.600 473.640 ;
        RECT 3.990 470.240 1196.000 472.240 ;
        RECT 3.990 468.840 1195.600 470.240 ;
        RECT 3.990 466.840 1196.000 468.840 ;
        RECT 3.990 465.440 1195.600 466.840 ;
        RECT 3.990 463.440 1196.000 465.440 ;
        RECT 3.990 462.040 1195.600 463.440 ;
        RECT 3.990 460.040 1196.000 462.040 ;
        RECT 3.990 458.640 1195.600 460.040 ;
        RECT 3.990 456.640 1196.000 458.640 ;
        RECT 3.990 455.240 1195.600 456.640 ;
        RECT 3.990 453.240 1196.000 455.240 ;
        RECT 3.990 451.840 1195.600 453.240 ;
        RECT 3.990 449.840 1196.000 451.840 ;
        RECT 3.990 448.440 1195.600 449.840 ;
        RECT 3.990 446.440 1196.000 448.440 ;
        RECT 3.990 445.040 1195.600 446.440 ;
        RECT 3.990 443.040 1196.000 445.040 ;
        RECT 3.990 441.640 1195.600 443.040 ;
        RECT 3.990 439.640 1196.000 441.640 ;
        RECT 3.990 438.240 1195.600 439.640 ;
        RECT 3.990 10.715 1196.000 438.240 ;
      LAYER met4 ;
        RECT 749.175 472.095 788.640 1170.105 ;
        RECT 791.040 472.095 791.940 1170.105 ;
        RECT 794.340 472.095 942.240 1170.105 ;
        RECT 944.640 472.095 945.540 1170.105 ;
        RECT 947.940 472.095 1095.840 1170.105 ;
        RECT 1098.240 472.095 1099.140 1170.105 ;
        RECT 1101.540 472.095 1110.145 1170.105 ;
  END
END des_core
END LIBRARY

